module gpio_top_apb(
  input         clock,
  input         reset,
  input  [31:0] in_paddr,
  input         in_psel,
  input         in_penable,
  input  [2:0]  in_pprot,
  input         in_pwrite,
  input  [31:0] in_pwdata,
  input  [3:0]  in_pstrb,
  output        in_pready,
  output [31:0] in_prdata,
  output        in_pslverr,

  output [15:0] gpio_out,
  input  [15:0] gpio_in,
  output [7:0]  gpio_seg_0,
  output [7:0]  gpio_seg_1,
  output [7:0]  gpio_seg_2,
  output [7:0]  gpio_seg_3,
  output [7:0]  gpio_seg_4,
  output [7:0]  gpio_seg_5,
  output [7:0]  gpio_seg_6,
  output [7:0]  gpio_seg_7
);

  reg [15:0] gpio_led;
  reg [31:0] gpio_seg;
  always @(posedge clock) begin
    if (reset) begin
      gpio_led <= 16'h0;
      gpio_seg <= 32'h0;
    end else if (in_penable && in_pwrite) begin
      if (in_paddr == 32'h10002000) begin
        gpio_led <= in_pwdata[15:0];
      end else if (in_paddr == 32'h10002008) begin
        gpio_seg <= in_pwdata;
      end
    end
  end
      
  assign gpio_out = gpio_led;
  assign in_pready = 1'b1;
  assign in_pslverr = 1'b0;
  assign in_prdata = {16'h0, gpio_in};

  assign gpio_seg_0 = {8{gpio_seg[3:0] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[3:0] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[3:0] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[3:0] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[3:0] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[3:0] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[3:0] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[3:0] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[3:0] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[3:0] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[3:0] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[3:0] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[3:0] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[3:0] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[3:0] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[3:0] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_1 = {8{gpio_seg[7:4] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[7:4] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[7:4] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[7:4] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[7:4] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[7:4] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[7:4] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[7:4] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[7:4] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[7:4] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[7:4] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[7:4] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[7:4] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[7:4] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[7:4] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[7:4] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_2 = {8{gpio_seg[11:8] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[11:8] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[11:8] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[11:8] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[11:8] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[11:8] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[11:8] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[11:8] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[11:8] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[11:8] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[11:8] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[11:8] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[11:8] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[11:8] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[11:8] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[11:8] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_3 = {8{gpio_seg[15:12] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[15:12] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[15:12] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[15:12] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[15:12] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[15:12] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[15:12] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[15:12] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[15:12] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[15:12] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[15:12] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[15:12] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[15:12] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[15:12] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[15:12] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[15:12] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_4 = {8{gpio_seg[19:16] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[19:16] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[19:16] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[19:16] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[19:16] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[19:16] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[19:16] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[19:16] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[19:16] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[19:16] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[19:16] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[19:16] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[19:16] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[19:16] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[19:16] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[19:16] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_5 = {8{gpio_seg[23:20] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[23:20] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[23:20] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[23:20] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[23:20] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[23:20] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[23:20] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[23:20] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[23:20] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[23:20] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[23:20] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[23:20] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[23:20] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[23:20] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[23:20] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[23:20] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_6 = {8{gpio_seg[27:24] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[27:24] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[27:24] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[27:24] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[27:24] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[27:24] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[27:24] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[27:24] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[27:24] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[27:24] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[27:24] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[27:24] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[27:24] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[27:24] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[27:24] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[27:24] == 4'b1111}} & 8'b01110001;

  assign gpio_seg_7 = {8{gpio_seg[31:28] == 4'b0000}} & 8'b00000011 |
                      {8{gpio_seg[31:28] == 4'b0001}} & 8'b10011111 |
                      {8{gpio_seg[31:28] == 4'b0010}} & 8'b00100101 |
                      {8{gpio_seg[31:28] == 4'b0011}} & 8'b00001101 |
                      {8{gpio_seg[31:28] == 4'b0100}} & 8'b10011001 |
                      {8{gpio_seg[31:28] == 4'b0101}} & 8'b01001001 |
                      {8{gpio_seg[31:28] == 4'b0110}} & 8'b01000001 |
                      {8{gpio_seg[31:28] == 4'b0111}} & 8'b00011111 |
                      {8{gpio_seg[31:28] == 4'b1000}} & 8'b00000001 |
                      {8{gpio_seg[31:28] == 4'b1001}} & 8'b00001001 |
                      {8{gpio_seg[31:28] == 4'b1010}} & 8'b00010001 |
                      {8{gpio_seg[31:28] == 4'b1011}} & 8'b11000001 |
                      {8{gpio_seg[31:28] == 4'b1100}} & 8'b01100011 |
                      {8{gpio_seg[31:28] == 4'b1101}} & 8'b10000101 |
                      {8{gpio_seg[31:28] == 4'b1110}} & 8'b01100001 |
                      {8{gpio_seg[31:28] == 4'b1111}} & 8'b01110001;
endmodule
