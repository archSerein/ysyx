module execute (
    input                               clk_i,
    input                               rst_i,
    input                               mem_valid_i,
    input  [`MEM_EXECUTE_BUS_WIDTH-1:0] mem_execute_bus_i,
    output [`EXECUTE_WB_BUS_WIDTH-1:0]  execute_wb_bus_o,
    output                              valid_o
);


endmodule